// Package file , contains all .sv files

`include "message_sender.sv";
`include "message_receiver.sv";
`include "message_test.sv";

